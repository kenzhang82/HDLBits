module counter1to12
(
	input clk,
	input reset,
	input enable,
	output [3:0] Q,
	output c_enable,
	output c_load,
	output [3:0] c_d
);

  
	count4 count4_inst
	(
		.clk(clk),
		.enable(c_enable),
		.load(c_load),
		.d(c_d),
		.Q(Q)
	);

  assign c_enable = enable;
  assign c_load = reset || (Q == 4'd12);
  assign c_d = 1;

endmodule
module shift4 
(
  input clk,
  input areset,
  input load,
  input ena,
  input [3:0] data,
  output reg [3:0] q 
);
  
  // TODO

endmodule
module countslow
(
	input clk,
	input slowena,
	input reset,
	output [3:0] q
);

	always @(posedge clk) begin
		if (reset) begin
			q <= 0;
		end
		else begin
			if (slowena) begin
				if (q < 4'd9) begin
					q <= q + 1;
				end
				else begin
					q <= 0;
				end
			end
		end
	end

endmodule
module wire
(
	input in,
	output out
);

	assign out = in;

endmodule